library IEEE;
use IEEE.STD_LOGIC_1164.all;
--library xil_defaultlib;


package wb_switch_pkg is

	constant MAX_OFFSETS		: natural := 8;

	type offsets_arr_t is array (0 to MAX_OFFSETS) of natural;
	end wb_switch_pkg;

package body wb_switch_pkg is
end wb_switch_pkg;
